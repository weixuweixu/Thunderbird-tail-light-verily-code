magic
tech scmos
timestamp 1520029804
<< metal1 >>
rect 14 807 954 827
rect 38 783 930 803
rect 38 767 930 773
rect 266 743 276 746
rect 124 733 132 736
rect 250 726 253 735
rect 284 733 293 736
rect 130 723 140 726
rect 180 723 189 726
rect 236 723 253 726
rect 260 723 277 726
rect 308 723 324 726
rect 338 723 348 726
rect 578 723 588 726
rect 338 715 341 723
rect 14 667 954 673
rect 178 633 188 636
rect 196 623 205 626
rect 580 623 588 626
rect 660 623 708 626
rect 810 616 813 625
rect 108 613 125 616
rect 164 613 180 616
rect 274 613 284 616
rect 314 606 317 614
rect 340 613 349 616
rect 436 613 461 616
rect 514 606 517 614
rect 548 613 564 616
rect 730 613 740 616
rect 746 613 756 616
rect 770 613 788 616
rect 802 613 813 616
rect 834 613 844 616
rect 308 603 317 606
rect 338 603 396 606
rect 410 603 420 606
rect 444 603 517 606
rect 530 603 540 606
rect 730 605 733 613
rect 748 603 757 606
rect 764 603 780 606
rect 802 605 805 613
rect 834 605 837 613
rect 466 593 492 596
rect 530 595 533 603
rect 38 567 930 573
rect 308 533 317 536
rect 348 533 357 536
rect 370 533 388 536
rect 474 533 484 536
rect 108 523 125 526
rect 290 523 301 526
rect 370 525 373 533
rect 530 526 533 535
rect 708 533 717 536
rect 530 523 549 526
rect 612 523 636 526
rect 652 523 685 526
rect 714 525 717 533
rect 738 533 748 536
rect 738 525 741 533
rect 778 526 781 535
rect 812 533 821 536
rect 778 523 789 526
rect 810 523 820 526
rect 290 515 293 523
rect 786 515 789 523
rect 14 467 954 473
rect 620 433 629 436
rect 90 416 93 425
rect 554 416 557 425
rect 604 423 612 426
rect 84 413 93 416
rect 148 413 157 416
rect 308 413 324 416
rect 338 413 356 416
rect 524 413 532 416
rect 546 413 557 416
rect 564 413 588 416
rect 554 406 557 413
rect 66 403 76 406
rect 282 403 300 406
rect 466 403 516 406
rect 546 403 557 406
rect 674 403 764 406
rect 546 395 549 403
rect 706 393 756 396
rect 38 367 930 373
rect 474 343 508 346
rect 690 336 693 345
rect 404 333 413 336
rect 420 333 429 336
rect 524 333 533 336
rect 604 333 621 336
rect 642 333 652 336
rect 666 333 676 336
rect 690 333 700 336
rect 466 323 508 326
rect 548 323 557 326
rect 618 325 621 333
rect 722 326 725 335
rect 778 326 781 335
rect 644 323 653 326
rect 722 323 732 326
rect 738 323 748 326
rect 772 323 781 326
rect 826 326 829 345
rect 826 323 836 326
rect 554 316 557 323
rect 554 313 564 316
rect 14 267 954 273
rect 666 216 669 225
rect 754 216 757 225
rect 114 206 117 214
rect 194 206 197 214
rect 268 213 285 216
rect 324 213 333 216
rect 340 213 349 216
rect 370 213 381 216
rect 114 203 124 206
rect 154 203 164 206
rect 194 203 204 206
rect 330 205 333 213
rect 378 205 381 213
rect 402 213 412 216
rect 498 213 516 216
rect 522 213 540 216
rect 580 213 597 216
rect 636 213 645 216
rect 652 213 669 216
rect 684 213 693 216
rect 754 213 772 216
rect 402 205 405 213
rect 490 203 508 206
rect 642 205 645 213
rect 658 203 668 206
rect 692 203 732 206
rect 756 203 765 206
rect 38 167 930 173
rect 148 133 156 136
rect 202 126 205 135
rect 402 126 405 135
rect 418 133 428 136
rect 452 133 484 136
rect 508 133 517 136
rect 530 126 533 135
rect 770 126 773 135
rect 786 133 796 136
rect 116 123 133 126
rect 178 123 205 126
rect 226 123 244 126
rect 340 123 357 126
rect 396 123 405 126
rect 412 123 429 126
rect 444 123 461 126
rect 506 123 524 126
rect 530 123 540 126
rect 578 123 596 126
rect 708 123 725 126
rect 764 123 773 126
rect 780 123 797 126
rect 812 123 836 126
rect 178 115 181 123
rect 226 115 229 123
rect 426 115 429 123
rect 506 115 509 123
rect 794 115 797 123
rect 14 67 954 73
rect 38 37 930 57
rect 14 13 954 33
<< metal2 >>
rect 14 13 34 827
rect 38 37 58 803
rect 114 743 117 840
rect 82 533 85 616
rect 122 583 125 616
rect 130 613 133 756
rect 154 733 157 756
rect 250 743 269 746
rect 250 733 253 743
rect 290 733 293 746
rect 154 566 157 586
rect 170 576 173 626
rect 150 563 157 566
rect 162 573 173 576
rect 66 393 69 406
rect 74 353 85 356
rect 82 333 85 353
rect 98 276 101 416
rect 106 403 109 516
rect 122 503 125 526
rect 150 516 153 563
rect 162 523 165 573
rect 178 566 181 636
rect 186 613 189 726
rect 170 563 181 566
rect 170 523 173 563
rect 150 513 157 516
rect 202 513 205 626
rect 154 426 157 513
rect 154 423 165 426
rect 122 353 125 406
rect 154 396 157 416
rect 150 393 157 396
rect 106 306 109 326
rect 150 316 153 393
rect 162 323 165 423
rect 178 333 181 356
rect 202 353 205 506
rect 226 503 229 526
rect 250 476 253 546
rect 266 533 269 626
rect 274 613 277 726
rect 290 713 293 726
rect 298 626 301 736
rect 314 733 317 746
rect 338 723 341 736
rect 402 723 405 746
rect 426 733 429 756
rect 442 733 445 746
rect 298 623 309 626
rect 274 593 277 606
rect 282 586 285 616
rect 290 603 293 616
rect 298 603 301 616
rect 306 593 309 623
rect 282 583 301 586
rect 290 533 293 576
rect 242 473 253 476
rect 242 376 245 473
rect 242 373 249 376
rect 150 313 157 316
rect 106 303 117 306
rect 90 273 101 276
rect 90 216 93 273
rect 114 246 117 303
rect 106 243 117 246
rect 90 213 101 216
rect 98 183 101 213
rect 106 203 109 243
rect 122 196 125 226
rect 138 203 141 216
rect 122 193 141 196
rect 82 133 85 146
rect 130 133 133 156
rect 130 113 133 126
rect 138 123 141 193
rect 146 146 149 206
rect 154 203 157 313
rect 202 266 205 326
rect 246 316 249 373
rect 258 323 261 506
rect 274 436 277 526
rect 298 523 301 583
rect 314 533 317 596
rect 322 533 325 716
rect 338 663 341 716
rect 442 713 445 726
rect 330 583 333 606
rect 314 513 317 526
rect 330 523 333 546
rect 338 516 341 606
rect 346 573 349 616
rect 354 543 357 586
rect 338 513 349 516
rect 354 486 357 536
rect 362 513 365 546
rect 370 533 373 556
rect 378 523 381 666
rect 386 613 389 626
rect 402 593 405 616
rect 426 613 429 706
rect 458 613 461 726
rect 466 703 469 736
rect 530 723 533 736
rect 562 733 565 840
rect 506 613 509 626
rect 402 536 405 586
rect 410 563 413 606
rect 402 533 421 536
rect 394 523 405 526
rect 346 483 357 486
rect 274 433 285 436
rect 282 323 285 433
rect 314 403 317 416
rect 322 413 325 426
rect 338 423 341 436
rect 330 413 341 416
rect 338 323 341 406
rect 346 403 349 483
rect 362 423 365 476
rect 370 413 373 426
rect 378 413 381 436
rect 386 366 389 426
rect 394 423 397 516
rect 410 433 413 526
rect 418 473 421 533
rect 426 516 429 546
rect 426 513 437 516
rect 426 453 429 513
rect 442 426 445 566
rect 450 503 453 606
rect 466 593 469 606
rect 522 563 525 606
rect 458 433 461 516
rect 394 413 405 416
rect 386 363 405 366
rect 418 363 421 426
rect 442 423 453 426
rect 246 313 253 316
rect 186 263 205 266
rect 154 183 157 196
rect 146 143 157 146
rect 146 106 149 136
rect 138 103 149 106
rect 138 86 141 103
rect 130 83 141 86
rect 130 16 133 83
rect 130 13 141 16
rect 138 0 141 13
rect 154 0 157 143
rect 162 126 165 206
rect 170 186 173 216
rect 186 203 189 263
rect 250 256 253 313
rect 242 253 253 256
rect 178 193 189 196
rect 170 183 181 186
rect 186 183 189 193
rect 178 133 181 183
rect 186 133 189 156
rect 162 123 181 126
rect 178 0 181 123
rect 194 113 197 146
rect 202 136 205 226
rect 218 143 221 216
rect 226 146 229 206
rect 242 183 245 253
rect 282 193 285 216
rect 226 143 245 146
rect 202 133 229 136
rect 202 123 213 126
rect 234 103 237 136
rect 242 123 245 143
rect 314 133 317 236
rect 362 233 365 336
rect 378 333 381 346
rect 386 323 389 356
rect 402 313 405 363
rect 426 356 429 416
rect 434 413 445 416
rect 410 333 413 356
rect 418 353 429 356
rect 418 326 421 353
rect 434 346 437 406
rect 450 403 453 423
rect 426 343 437 346
rect 426 333 437 336
rect 410 323 421 326
rect 346 223 373 226
rect 346 213 365 216
rect 370 213 373 223
rect 378 206 381 226
rect 330 166 333 206
rect 346 193 349 206
rect 370 203 381 206
rect 394 183 397 216
rect 410 213 413 323
rect 418 296 421 316
rect 434 313 437 333
rect 442 323 445 366
rect 466 333 469 406
rect 474 403 477 536
rect 514 513 517 526
rect 530 516 533 616
rect 554 603 557 626
rect 578 603 581 726
rect 594 633 597 736
rect 610 733 613 756
rect 706 733 709 756
rect 802 733 805 756
rect 538 533 549 536
rect 554 533 557 546
rect 562 526 565 566
rect 530 513 541 516
rect 482 436 485 456
rect 482 433 493 436
rect 490 386 493 433
rect 530 396 533 416
rect 538 406 541 513
rect 546 496 549 526
rect 554 523 565 526
rect 554 513 557 523
rect 570 513 573 576
rect 578 506 581 536
rect 586 533 589 626
rect 602 533 605 616
rect 610 606 613 626
rect 626 623 637 626
rect 610 603 621 606
rect 626 603 629 616
rect 618 573 621 603
rect 642 573 645 616
rect 650 583 653 636
rect 586 523 597 526
rect 570 503 581 506
rect 610 503 613 526
rect 618 513 621 536
rect 626 533 629 566
rect 642 533 645 546
rect 546 493 557 496
rect 554 436 557 493
rect 546 433 557 436
rect 546 413 549 433
rect 538 403 549 406
rect 530 393 541 396
rect 482 383 493 386
rect 474 343 477 356
rect 442 313 461 316
rect 418 293 425 296
rect 422 226 425 293
rect 418 223 425 226
rect 418 203 421 223
rect 434 203 437 216
rect 442 203 445 313
rect 466 306 469 326
rect 482 313 485 383
rect 450 303 469 306
rect 434 183 437 196
rect 330 163 341 166
rect 338 86 341 163
rect 354 123 357 146
rect 418 133 421 146
rect 330 83 341 86
rect 330 0 333 83
rect 402 0 405 126
rect 418 113 421 126
rect 450 123 453 216
rect 458 123 461 206
rect 490 203 493 366
rect 522 326 525 336
rect 530 333 533 346
rect 522 323 533 326
rect 522 223 525 316
rect 538 313 541 393
rect 570 356 573 503
rect 578 393 581 406
rect 602 403 605 426
rect 610 413 613 426
rect 618 406 621 436
rect 626 433 629 526
rect 634 423 637 526
rect 610 403 621 406
rect 570 353 581 356
rect 546 313 549 326
rect 554 323 557 336
rect 562 333 565 346
rect 578 323 581 353
rect 586 333 589 356
rect 594 323 597 376
rect 610 343 613 403
rect 626 393 629 416
rect 626 323 629 386
rect 634 336 637 416
rect 658 383 661 626
rect 706 623 709 636
rect 706 603 709 616
rect 682 533 685 556
rect 722 533 725 616
rect 730 613 733 726
rect 786 626 789 726
rect 786 623 797 626
rect 682 503 685 526
rect 690 493 693 526
rect 642 343 661 346
rect 634 333 645 336
rect 650 303 653 326
rect 658 323 661 343
rect 666 333 669 346
rect 674 326 677 406
rect 706 393 709 516
rect 738 383 741 586
rect 746 566 749 616
rect 770 606 773 616
rect 754 603 773 606
rect 770 583 773 596
rect 746 563 757 566
rect 754 523 757 563
rect 762 423 765 536
rect 786 533 789 616
rect 794 583 797 623
rect 802 596 805 716
rect 826 676 829 726
rect 882 713 885 726
rect 810 673 829 676
rect 810 603 813 673
rect 826 613 829 636
rect 802 593 813 596
rect 770 493 773 526
rect 802 523 805 536
rect 786 503 789 516
rect 698 333 701 366
rect 666 323 677 326
rect 490 123 493 196
rect 498 183 501 216
rect 522 193 525 216
rect 530 183 533 206
rect 554 183 557 236
rect 594 193 597 216
rect 658 213 661 226
rect 690 213 693 326
rect 714 323 717 346
rect 738 333 741 356
rect 746 343 749 366
rect 698 303 701 316
rect 738 306 741 326
rect 730 303 741 306
rect 730 236 733 303
rect 730 233 741 236
rect 514 133 517 146
rect 514 113 517 126
rect 538 0 541 126
rect 578 123 581 146
rect 618 133 621 186
rect 642 156 645 206
rect 658 193 661 206
rect 642 153 653 156
rect 650 106 653 153
rect 682 133 685 146
rect 698 123 701 216
rect 738 213 741 233
rect 754 183 757 376
rect 762 333 765 356
rect 770 336 773 436
rect 810 433 813 593
rect 834 556 837 606
rect 826 553 837 556
rect 818 533 821 546
rect 826 533 829 553
rect 834 513 837 526
rect 842 493 845 536
rect 850 456 853 606
rect 858 493 861 526
rect 866 516 869 546
rect 866 513 877 516
rect 850 453 857 456
rect 810 413 813 426
rect 786 373 789 406
rect 770 333 789 336
rect 794 333 805 336
rect 778 303 781 326
rect 786 313 789 333
rect 810 323 813 386
rect 818 316 821 336
rect 802 313 821 316
rect 762 213 765 226
rect 762 193 765 206
rect 778 203 781 226
rect 794 183 797 206
rect 818 193 821 216
rect 722 123 725 146
rect 786 133 789 146
rect 642 103 653 106
rect 642 0 645 103
rect 770 0 773 126
rect 786 113 789 126
rect 818 123 821 136
rect 826 133 829 366
rect 854 346 857 453
rect 874 436 877 513
rect 842 333 845 346
rect 850 343 857 346
rect 866 433 877 436
rect 850 303 853 343
rect 858 313 861 326
rect 866 303 869 433
rect 874 313 877 346
rect 874 213 877 226
rect 910 37 930 803
rect 934 13 954 827
<< metal3 >>
rect 273 772 406 777
rect 273 757 278 772
rect 129 752 278 757
rect 401 757 406 772
rect 513 762 590 767
rect 513 757 518 762
rect 401 752 518 757
rect 585 757 590 762
rect 585 752 806 757
rect 289 742 318 747
rect 401 742 446 747
rect 529 732 598 737
rect 337 722 446 727
rect 289 712 326 717
rect 801 712 886 717
rect 425 702 470 707
rect 337 662 382 667
rect 289 632 366 637
rect 289 627 294 632
rect 265 622 294 627
rect 361 627 366 632
rect 409 632 486 637
rect 705 632 830 637
rect 409 627 414 632
rect 361 622 414 627
rect 481 627 486 632
rect 481 622 662 627
rect 81 612 134 617
rect 185 612 294 617
rect 401 612 534 617
rect 705 612 734 617
rect 297 602 750 607
rect 273 592 342 597
rect 721 592 838 597
rect 121 582 270 587
rect 329 582 406 587
rect 649 582 742 587
rect 769 582 854 587
rect 289 572 350 577
rect 569 572 646 577
rect 313 562 446 567
rect 521 562 566 567
rect 625 562 662 567
rect 297 552 374 557
rect 681 552 814 557
rect 81 542 254 547
rect 329 542 366 547
rect 377 542 430 547
rect 553 542 646 547
rect 817 542 870 547
rect 537 532 614 537
rect 753 532 806 537
rect 609 527 614 532
rect 401 522 590 527
rect 609 522 630 527
rect 649 517 814 522
rect 105 512 206 517
rect 273 512 342 517
rect 361 512 398 517
rect 513 512 574 517
rect 617 512 654 517
rect 809 512 838 517
rect 337 507 342 512
rect 121 502 206 507
rect 225 502 262 507
rect 337 502 414 507
rect 577 502 614 507
rect 681 502 790 507
rect 633 492 694 497
rect 705 492 862 497
rect 361 472 422 477
rect 425 452 486 457
rect 337 432 462 437
rect 769 432 814 437
rect 321 422 374 427
rect 481 422 606 427
rect 761 422 814 427
rect 481 417 486 422
rect 313 412 334 417
rect 377 412 486 417
rect 609 412 638 417
rect 0 402 70 407
rect 433 402 550 407
rect 65 392 70 402
rect 537 392 630 397
rect 625 382 662 387
rect 737 382 814 387
rect 465 372 598 377
rect 753 372 790 377
rect 241 362 366 367
rect 417 362 494 367
rect 697 362 830 367
rect 241 357 246 362
rect 0 352 182 357
rect 201 352 246 357
rect 361 357 366 362
rect 361 352 390 357
rect 409 352 478 357
rect 513 352 614 357
rect 689 352 766 357
rect 513 347 518 352
rect 689 347 694 352
rect 257 342 286 347
rect 281 337 286 342
rect 353 342 518 347
rect 529 342 694 347
rect 713 342 878 347
rect 353 337 358 342
rect 281 332 358 337
rect 385 332 470 337
rect 521 332 654 337
rect 649 327 654 332
rect 761 332 798 337
rect 761 327 766 332
rect 553 322 630 327
rect 649 322 766 327
rect 417 312 486 317
rect 521 312 550 317
rect 785 312 862 317
rect 649 302 702 307
rect 777 302 854 307
rect 385 242 462 247
rect 385 237 390 242
rect 313 232 390 237
rect 457 237 462 242
rect 457 232 558 237
rect 777 222 902 227
rect 897 217 902 222
rect 377 212 446 217
rect 657 212 766 217
rect 897 212 968 217
rect 137 202 166 207
rect 433 202 462 207
rect 281 192 350 197
rect 489 192 526 197
rect 593 192 662 197
rect 761 192 822 197
rect 97 182 190 187
rect 241 182 318 187
rect 393 182 534 187
rect 553 182 798 187
rect 129 152 190 157
rect 81 142 142 147
rect 193 142 222 147
rect 353 142 422 147
rect 513 142 582 147
rect 617 142 686 147
rect 721 142 790 147
rect 137 127 142 137
rect 137 122 206 127
rect 417 122 542 127
rect 537 117 542 122
rect 673 122 822 127
rect 673 117 678 122
rect 129 112 198 117
rect 537 112 678 117
rect 177 102 238 107
use turn_VIA1  turn_VIA1_0
timestamp 1520029804
transform 1 0 24 0 1 817
box -10 -10 10 10
use turn_VIA1  turn_VIA1_1
timestamp 1520029804
transform 1 0 944 0 1 817
box -10 -10 10 10
use turn_VIA1  turn_VIA1_2
timestamp 1520029804
transform 1 0 48 0 1 793
box -10 -10 10 10
use turn_VIA1  turn_VIA1_3
timestamp 1520029804
transform 1 0 920 0 1 793
box -10 -10 10 10
use turn_VIA0  turn_VIA0_0
timestamp 1520029804
transform 1 0 48 0 1 770
box -10 -3 10 3
use M2_M1  M2_M1_0
timestamp 1520029804
transform 1 0 116 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1520029804
transform 1 0 132 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_14
timestamp 1520029804
transform 1 0 132 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_1
timestamp 1520029804
transform 1 0 156 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_2
timestamp 1520029804
transform 1 0 156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1520029804
transform 1 0 188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1520029804
transform 1 0 252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1520029804
transform 1 0 268 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1520029804
transform 1 0 276 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_6
timestamp 1520029804
transform 1 0 292 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1520029804
transform 1 0 316 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4
timestamp 1520029804
transform 1 0 292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1520029804
transform 1 0 300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1520029804
transform 1 0 316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1520029804
transform 1 0 292 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_2
timestamp 1520029804
transform 1 0 428 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1520029804
transform 1 0 404 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1520029804
transform 1 0 444 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_7
timestamp 1520029804
transform 1 0 340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1520029804
transform 1 0 428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1520029804
transform 1 0 444 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_13
timestamp 1520029804
transform 1 0 340 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_18
timestamp 1520029804
transform 1 0 404 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_15
timestamp 1520029804
transform 1 0 292 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1520029804
transform 1 0 324 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_26
timestamp 1520029804
transform 1 0 340 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_14
timestamp 1520029804
transform 1 0 444 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1520029804
transform 1 0 468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1520029804
transform 1 0 460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1520029804
transform 1 0 444 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_19
timestamp 1520029804
transform 1 0 428 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1520029804
transform 1 0 468 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1520029804
transform 1 0 612 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1520029804
transform 1 0 532 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1520029804
transform 1 0 564 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1520029804
transform 1 0 596 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1520029804
transform 1 0 612 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1520029804
transform 1 0 532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1520029804
transform 1 0 580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_4
timestamp 1520029804
transform 1 0 708 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_12
timestamp 1520029804
transform 1 0 708 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_5
timestamp 1520029804
transform 1 0 804 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1520029804
transform 1 0 804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1520029804
transform 1 0 732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1520029804
transform 1 0 788 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1520029804
transform 1 0 828 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1520029804
transform 1 0 884 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_17
timestamp 1520029804
transform 1 0 804 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1520029804
transform 1 0 884 0 1 715
box -3 -3 3 3
use turn_VIA0  turn_VIA0_1
timestamp 1520029804
transform 1 0 920 0 1 770
box -10 -3 10 3
use turn_VIA0  turn_VIA0_2
timestamp 1520029804
transform 1 0 24 0 1 670
box -10 -3 10 3
use FILL  FILL_0
timestamp 1520029804
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_1
timestamp 1520029804
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_2
timestamp 1520029804
transform 1 0 88 0 -1 770
box -8 -3 16 105
use FILL  FILL_3
timestamp 1520029804
transform 1 0 96 0 -1 770
box -8 -3 16 105
use FILL  FILL_4
timestamp 1520029804
transform 1 0 104 0 -1 770
box -8 -3 16 105
use INVX1  INVX1_0
timestamp 1520029804
transform 1 0 112 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_0
timestamp 1520029804
transform 1 0 128 0 -1 770
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_0
timestamp 1520029804
transform 1 0 144 0 -1 770
box -8 -3 104 105
use FILL  FILL_5
timestamp 1520029804
transform 1 0 240 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_1
timestamp 1520029804
transform 1 0 248 0 -1 770
box -9 -3 26 105
use FILL  FILL_6
timestamp 1520029804
transform 1 0 264 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1520029804
transform 1 0 272 0 -1 770
box -8 -3 32 105
use INVX2  INVX2_2
timestamp 1520029804
transform 1 0 296 0 -1 770
box -9 -3 26 105
use OAI21X1  OAI21X1_0
timestamp 1520029804
transform 1 0 312 0 -1 770
box -8 -3 34 105
use DFFPOSX1  DFFPOSX1_1
timestamp 1520029804
transform -1 0 440 0 -1 770
box -8 -3 104 105
use OAI21X1  OAI21X1_1
timestamp 1520029804
transform -1 0 472 0 -1 770
box -8 -3 34 105
use FILL  FILL_7
timestamp 1520029804
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_8
timestamp 1520029804
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_9
timestamp 1520029804
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_10
timestamp 1520029804
transform 1 0 496 0 -1 770
box -8 -3 16 105
use FILL  FILL_11
timestamp 1520029804
transform 1 0 504 0 -1 770
box -8 -3 16 105
use FILL  FILL_12
timestamp 1520029804
transform 1 0 512 0 -1 770
box -8 -3 16 105
use FILL  FILL_13
timestamp 1520029804
transform 1 0 520 0 -1 770
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_2
timestamp 1520029804
transform -1 0 624 0 -1 770
box -8 -3 104 105
use FILL  FILL_14
timestamp 1520029804
transform 1 0 624 0 -1 770
box -8 -3 16 105
use FILL  FILL_15
timestamp 1520029804
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_16
timestamp 1520029804
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_17
timestamp 1520029804
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_18
timestamp 1520029804
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_19
timestamp 1520029804
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_20
timestamp 1520029804
transform 1 0 672 0 -1 770
box -8 -3 16 105
use FILL  FILL_21
timestamp 1520029804
transform 1 0 680 0 -1 770
box -8 -3 16 105
use FILL  FILL_22
timestamp 1520029804
transform 1 0 688 0 -1 770
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_3
timestamp 1520029804
transform 1 0 696 0 -1 770
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_4
timestamp 1520029804
transform 1 0 792 0 -1 770
box -8 -3 104 105
use FILL  FILL_23
timestamp 1520029804
transform 1 0 888 0 -1 770
box -8 -3 16 105
use turn_VIA0  turn_VIA0_3
timestamp 1520029804
transform 1 0 944 0 1 670
box -10 -3 10 3
use M2_M1  M2_M1_28
timestamp 1520029804
transform 1 0 180 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1520029804
transform 1 0 172 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_32
timestamp 1520029804
transform 1 0 84 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1520029804
transform 1 0 124 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_33
timestamp 1520029804
transform 1 0 132 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_54
timestamp 1520029804
transform 1 0 84 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_50
timestamp 1520029804
transform 1 0 124 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1520029804
transform 1 0 156 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1520029804
transform 1 0 188 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_32
timestamp 1520029804
transform 1 0 204 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_25
timestamp 1520029804
transform 1 0 268 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_38
timestamp 1520029804
transform 1 0 276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1520029804
transform 1 0 284 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_35
timestamp 1520029804
transform 1 0 292 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_40
timestamp 1520029804
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1520029804
transform 1 0 276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1520029804
transform 1 0 292 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_40
timestamp 1520029804
transform 1 0 300 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1520029804
transform 1 0 276 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1520029804
transform 1 0 268 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1520029804
transform 1 0 340 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1520029804
transform 1 0 324 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_41
timestamp 1520029804
transform 1 0 348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1520029804
transform 1 0 332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1520029804
transform 1 0 340 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_46
timestamp 1520029804
transform 1 0 308 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_71
timestamp 1520029804
transform 1 0 316 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_47
timestamp 1520029804
transform 1 0 340 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1520029804
transform 1 0 332 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1520029804
transform 1 0 356 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1520029804
transform 1 0 380 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1520029804
transform 1 0 388 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_42
timestamp 1520029804
transform 1 0 388 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_36
timestamp 1520029804
transform 1 0 404 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_59
timestamp 1520029804
transform 1 0 412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1520029804
transform 1 0 404 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_55
timestamp 1520029804
transform 1 0 404 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1520029804
transform 1 0 428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1520029804
transform 1 0 452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1520029804
transform 1 0 460 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1520029804
transform 1 0 468 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_73
timestamp 1520029804
transform 1 0 468 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_27
timestamp 1520029804
transform 1 0 508 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_45
timestamp 1520029804
transform 1 0 508 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_28
timestamp 1520029804
transform 1 0 556 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1520029804
transform 1 0 532 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_61
timestamp 1520029804
transform 1 0 524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1520029804
transform 1 0 532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1520029804
transform 1 0 556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1520029804
transform 1 0 596 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_29
timestamp 1520029804
transform 1 0 588 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_30
timestamp 1520029804
transform 1 0 652 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1520029804
transform 1 0 612 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1520029804
transform 1 0 604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1520029804
transform 1 0 580 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_30
timestamp 1520029804
transform 1 0 628 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_34
timestamp 1520029804
transform 1 0 636 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_31
timestamp 1520029804
transform 1 0 660 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_47
timestamp 1520029804
transform 1 0 628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1520029804
transform 1 0 644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1520029804
transform 1 0 620 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_43
timestamp 1520029804
transform 1 0 628 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1520029804
transform 1 0 652 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1520029804
transform 1 0 708 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_35
timestamp 1520029804
transform 1 0 708 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_38
timestamp 1520029804
transform 1 0 708 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_49
timestamp 1520029804
transform 1 0 724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1520029804
transform 1 0 708 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_39
timestamp 1520029804
transform 1 0 732 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_50
timestamp 1520029804
transform 1 0 748 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1520029804
transform 1 0 748 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_67
timestamp 1520029804
transform 1 0 756 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1520029804
transform 1 0 724 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1520029804
transform 1 0 740 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_36
timestamp 1520029804
transform 1 0 804 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1520029804
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1520029804
transform 1 0 788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1520029804
transform 1 0 772 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_58
timestamp 1520029804
transform 1 0 772 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1520029804
transform 1 0 796 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1520029804
transform 1 0 828 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_53
timestamp 1520029804
transform 1 0 828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1520029804
transform 1 0 812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1520029804
transform 1 0 836 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1520029804
transform 1 0 852 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1520029804
transform 1 0 836 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1520029804
transform 1 0 852 0 1 585
box -3 -3 3 3
use turn_VIA0  turn_VIA0_4
timestamp 1520029804
transform 1 0 48 0 1 570
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_5
timestamp 1520029804
transform 1 0 72 0 1 570
box -8 -3 104 105
use NAND3X1  NAND3X1_0
timestamp 1520029804
transform 1 0 168 0 1 570
box -8 -3 40 105
use FILL  FILL_24
timestamp 1520029804
transform 1 0 200 0 1 570
box -8 -3 16 105
use FILL  FILL_25
timestamp 1520029804
transform 1 0 208 0 1 570
box -8 -3 16 105
use FILL  FILL_26
timestamp 1520029804
transform 1 0 216 0 1 570
box -8 -3 16 105
use FILL  FILL_27
timestamp 1520029804
transform 1 0 224 0 1 570
box -8 -3 16 105
use FILL  FILL_28
timestamp 1520029804
transform 1 0 232 0 1 570
box -8 -3 16 105
use FILL  FILL_29
timestamp 1520029804
transform 1 0 240 0 1 570
box -8 -3 16 105
use FILL  FILL_30
timestamp 1520029804
transform 1 0 248 0 1 570
box -8 -3 16 105
use FILL  FILL_31
timestamp 1520029804
transform 1 0 256 0 1 570
box -8 -3 16 105
use FILL  FILL_32
timestamp 1520029804
transform 1 0 264 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_61
timestamp 1520029804
transform 1 0 292 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_0
timestamp 1520029804
transform 1 0 272 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_62
timestamp 1520029804
transform 1 0 348 0 1 575
box -3 -3 3 3
use AOI21X1  AOI21X1_0
timestamp 1520029804
transform -1 0 344 0 1 570
box -7 -3 39 105
use FILL  FILL_33
timestamp 1520029804
transform 1 0 344 0 1 570
box -8 -3 16 105
use FILL  FILL_34
timestamp 1520029804
transform 1 0 352 0 1 570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1520029804
transform 1 0 360 0 1 570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1520029804
transform 1 0 368 0 1 570
box -8 -3 16 105
use FILL  FILL_37
timestamp 1520029804
transform 1 0 376 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1520029804
transform -1 0 408 0 1 570
box -8 -3 32 105
use FILL  FILL_38
timestamp 1520029804
transform 1 0 408 0 1 570
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1520029804
transform 1 0 416 0 1 570
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1520029804
transform -1 0 448 0 1 570
box -9 -3 26 105
use FILL  FILL_39
timestamp 1520029804
transform 1 0 448 0 1 570
box -8 -3 16 105
use FILL  FILL_40
timestamp 1520029804
transform 1 0 456 0 1 570
box -8 -3 16 105
use FILL  FILL_41
timestamp 1520029804
transform 1 0 464 0 1 570
box -8 -3 16 105
use FILL  FILL_43
timestamp 1520029804
transform 1 0 472 0 1 570
box -8 -3 16 105
use FILL  FILL_45
timestamp 1520029804
transform 1 0 480 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1520029804
transform 1 0 488 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1520029804
transform -1 0 536 0 1 570
box -8 -3 32 105
use M3_M2  M3_M2_63
timestamp 1520029804
transform 1 0 572 0 1 575
box -3 -3 3 3
use INVX2  INVX2_6
timestamp 1520029804
transform 1 0 536 0 1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_4
timestamp 1520029804
transform 1 0 552 0 1 570
box -8 -3 34 105
use M3_M2  M3_M2_64
timestamp 1520029804
transform 1 0 620 0 1 575
box -3 -3 3 3
use NAND3X1  NAND3X1_2
timestamp 1520029804
transform -1 0 616 0 1 570
box -8 -3 40 105
use M3_M2  M3_M2_65
timestamp 1520029804
transform 1 0 644 0 1 575
box -3 -3 3 3
use INVX2  INVX2_7
timestamp 1520029804
transform 1 0 616 0 1 570
box -9 -3 26 105
use NAND3X1  NAND3X1_3
timestamp 1520029804
transform 1 0 632 0 1 570
box -8 -3 40 105
use FILL  FILL_46
timestamp 1520029804
transform 1 0 664 0 1 570
box -8 -3 16 105
use FILL  FILL_49
timestamp 1520029804
transform 1 0 672 0 1 570
box -8 -3 16 105
use FILL  FILL_51
timestamp 1520029804
transform 1 0 680 0 1 570
box -8 -3 16 105
use FILL  FILL_52
timestamp 1520029804
transform 1 0 688 0 1 570
box -8 -3 16 105
use FILL  FILL_53
timestamp 1520029804
transform 1 0 696 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1520029804
transform -1 0 736 0 1 570
box -8 -3 34 105
use INVX2  INVX2_11
timestamp 1520029804
transform -1 0 752 0 1 570
box -9 -3 26 105
use NOR2X1  NOR2X1_6
timestamp 1520029804
transform -1 0 776 0 1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_7
timestamp 1520029804
transform 1 0 776 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1520029804
transform -1 0 840 0 1 570
box -8 -3 34 105
use INVX2  INVX2_12
timestamp 1520029804
transform -1 0 856 0 1 570
box -9 -3 26 105
use FILL  FILL_54
timestamp 1520029804
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_55
timestamp 1520029804
transform 1 0 864 0 1 570
box -8 -3 16 105
use FILL  FILL_56
timestamp 1520029804
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_58
timestamp 1520029804
transform 1 0 880 0 1 570
box -8 -3 16 105
use FILL  FILL_60
timestamp 1520029804
transform 1 0 888 0 1 570
box -8 -3 16 105
use turn_VIA0  turn_VIA0_5
timestamp 1520029804
transform 1 0 920 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_77
timestamp 1520029804
transform 1 0 84 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_78
timestamp 1520029804
transform 1 0 84 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_78
timestamp 1520029804
transform 1 0 252 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_79
timestamp 1520029804
transform 1 0 252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1520029804
transform 1 0 268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1520029804
transform 1 0 124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1520029804
transform 1 0 164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1520029804
transform 1 0 172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1520029804
transform 1 0 228 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_93
timestamp 1520029804
transform 1 0 108 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1520029804
transform 1 0 124 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1520029804
transform 1 0 204 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1520029804
transform 1 0 316 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1520029804
transform 1 0 300 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_75
timestamp 1520029804
transform 1 0 300 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1520029804
transform 1 0 292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1520029804
transform 1 0 276 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_95
timestamp 1520029804
transform 1 0 276 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1520029804
transform 1 0 204 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1520029804
transform 1 0 228 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1520029804
transform 1 0 260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1520029804
transform 1 0 332 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_82
timestamp 1520029804
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1520029804
transform 1 0 324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1520029804
transform 1 0 300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1520029804
transform 1 0 316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1520029804
transform 1 0 332 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_96
timestamp 1520029804
transform 1 0 316 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1520029804
transform 1 0 372 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_76
timestamp 1520029804
transform 1 0 356 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_80
timestamp 1520029804
transform 1 0 364 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1520029804
transform 1 0 380 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1520029804
transform 1 0 412 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_84
timestamp 1520029804
transform 1 0 356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1520029804
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1520029804
transform 1 0 372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1520029804
transform 1 0 404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1520029804
transform 1 0 380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1520029804
transform 1 0 396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1520029804
transform 1 0 348 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_97
timestamp 1520029804
transform 1 0 364 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1520029804
transform 1 0 404 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_116
timestamp 1520029804
transform 1 0 412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1520029804
transform 1 0 420 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_98
timestamp 1520029804
transform 1 0 396 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1520029804
transform 1 0 412 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1520029804
transform 1 0 444 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1520029804
transform 1 0 428 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_88
timestamp 1520029804
transform 1 0 428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1520029804
transform 1 0 444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1520029804
transform 1 0 436 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1520029804
transform 1 0 460 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1520029804
transform 1 0 452 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1520029804
transform 1 0 476 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_69
timestamp 1520029804
transform 1 0 524 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1520029804
transform 1 0 540 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1520029804
transform 1 0 564 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1520029804
transform 1 0 556 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_90
timestamp 1520029804
transform 1 0 548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1520029804
transform 1 0 556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1520029804
transform 1 0 516 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1520029804
transform 1 0 516 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_120
timestamp 1520029804
transform 1 0 548 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_71
timestamp 1520029804
transform 1 0 628 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_92
timestamp 1520029804
transform 1 0 580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1520029804
transform 1 0 588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1520029804
transform 1 0 604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1520029804
transform 1 0 620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1520029804
transform 1 0 628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1520029804
transform 1 0 572 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_91
timestamp 1520029804
transform 1 0 588 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_122
timestamp 1520029804
transform 1 0 596 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1520029804
transform 1 0 612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1520029804
transform 1 0 556 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_100
timestamp 1520029804
transform 1 0 572 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1520029804
transform 1 0 628 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1520029804
transform 1 0 620 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1520029804
transform 1 0 580 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1520029804
transform 1 0 612 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1520029804
transform 1 0 644 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_97
timestamp 1520029804
transform 1 0 644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1520029804
transform 1 0 636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_112
timestamp 1520029804
transform 1 0 636 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1520029804
transform 1 0 660 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1520029804
transform 1 0 684 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_98
timestamp 1520029804
transform 1 0 684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1520029804
transform 1 0 684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1520029804
transform 1 0 692 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_110
timestamp 1520029804
transform 1 0 684 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_77
timestamp 1520029804
transform 1 0 740 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1520029804
transform 1 0 724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1520029804
transform 1 0 708 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_113
timestamp 1520029804
transform 1 0 692 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1520029804
transform 1 0 708 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1520029804
transform 1 0 756 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1520029804
transform 1 0 812 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1520029804
transform 1 0 820 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_100
timestamp 1520029804
transform 1 0 764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1520029804
transform 1 0 788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1520029804
transform 1 0 756 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1520029804
transform 1 0 772 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_89
timestamp 1520029804
transform 1 0 804 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_102
timestamp 1520029804
transform 1 0 820 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1520029804
transform 1 0 828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1520029804
transform 1 0 844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1520029804
transform 1 0 804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1520029804
transform 1 0 812 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1520029804
transform 1 0 836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1520029804
transform 1 0 852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1520029804
transform 1 0 860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1520029804
transform 1 0 788 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_111
timestamp 1520029804
transform 1 0 788 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1520029804
transform 1 0 772 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1520029804
transform 1 0 836 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1520029804
transform 1 0 868 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_105
timestamp 1520029804
transform 1 0 868 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_116
timestamp 1520029804
transform 1 0 844 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1520029804
transform 1 0 860 0 1 495
box -3 -3 3 3
use turn_VIA0  turn_VIA0_6
timestamp 1520029804
transform 1 0 24 0 1 470
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_6
timestamp 1520029804
transform 1 0 72 0 -1 570
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_7
timestamp 1520029804
transform -1 0 264 0 -1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_2
timestamp 1520029804
transform 1 0 264 0 -1 570
box -8 -3 34 105
use NOR2X1  NOR2X1_2
timestamp 1520029804
transform 1 0 296 0 -1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_3
timestamp 1520029804
transform 1 0 320 0 -1 570
box -8 -3 34 105
use M3_M2  M3_M2_118
timestamp 1520029804
transform 1 0 364 0 1 475
box -3 -3 3 3
use NOR2X1  NOR2X1_3
timestamp 1520029804
transform 1 0 352 0 -1 570
box -8 -3 32 105
use M3_M2  M3_M2_119
timestamp 1520029804
transform 1 0 420 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_0
timestamp 1520029804
transform 1 0 376 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_5
timestamp 1520029804
transform -1 0 432 0 -1 570
box -9 -3 26 105
use NAND3X1  NAND3X1_1
timestamp 1520029804
transform 1 0 432 0 -1 570
box -8 -3 40 105
use FILL  FILL_42
timestamp 1520029804
transform 1 0 464 0 -1 570
box -8 -3 16 105
use FILL  FILL_44
timestamp 1520029804
transform 1 0 472 0 -1 570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_0
timestamp 1520029804
transform 1 0 480 0 -1 570
box -8 -3 64 105
use INVX2  INVX2_8
timestamp 1520029804
transform -1 0 552 0 -1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_5
timestamp 1520029804
transform -1 0 584 0 -1 570
box -8 -3 34 105
use OAI22X1  OAI22X1_1
timestamp 1520029804
transform -1 0 624 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_9
timestamp 1520029804
transform 1 0 624 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1520029804
transform 1 0 640 0 -1 570
box -9 -3 26 105
use FILL  FILL_47
timestamp 1520029804
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_48
timestamp 1520029804
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_50
timestamp 1520029804
transform 1 0 672 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1520029804
transform 1 0 680 0 -1 570
box -8 -3 34 105
use AOI21X1  AOI21X1_1
timestamp 1520029804
transform 1 0 712 0 -1 570
box -7 -3 39 105
use OAI22X1  OAI22X1_2
timestamp 1520029804
transform -1 0 784 0 -1 570
box -8 -3 46 105
use OAI21X1  OAI21X1_10
timestamp 1520029804
transform -1 0 816 0 -1 570
box -8 -3 34 105
use AOI22X1  AOI22X1_1
timestamp 1520029804
transform 1 0 816 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_13
timestamp 1520029804
transform -1 0 872 0 -1 570
box -9 -3 26 105
use FILL  FILL_57
timestamp 1520029804
transform 1 0 872 0 -1 570
box -8 -3 16 105
use FILL  FILL_59
timestamp 1520029804
transform 1 0 880 0 -1 570
box -8 -3 16 105
use FILL  FILL_61
timestamp 1520029804
transform 1 0 888 0 -1 570
box -8 -3 16 105
use turn_VIA0  turn_VIA0_7
timestamp 1520029804
transform 1 0 944 0 1 470
box -10 -3 10 3
use M2_M1  M2_M1_167
timestamp 1520029804
transform 1 0 68 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_140
timestamp 1520029804
transform 1 0 68 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_152
timestamp 1520029804
transform 1 0 100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1520029804
transform 1 0 156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1520029804
transform 1 0 204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1520029804
transform 1 0 108 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1520029804
transform 1 0 124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1520029804
transform 1 0 284 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_122
timestamp 1520029804
transform 1 0 340 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1520029804
transform 1 0 324 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_145
timestamp 1520029804
transform 1 0 340 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_131
timestamp 1520029804
transform 1 0 316 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_155
timestamp 1520029804
transform 1 0 324 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_132
timestamp 1520029804
transform 1 0 332 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_156
timestamp 1520029804
transform 1 0 340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1520029804
transform 1 0 316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1520029804
transform 1 0 380 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1520029804
transform 1 0 364 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_127
timestamp 1520029804
transform 1 0 372 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1520029804
transform 1 0 428 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_142
timestamp 1520029804
transform 1 0 412 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1520029804
transform 1 0 388 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1520029804
transform 1 0 396 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1520029804
transform 1 0 340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1520029804
transform 1 0 348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1520029804
transform 1 0 372 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_133
timestamp 1520029804
transform 1 0 380 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1520029804
transform 1 0 396 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_149
timestamp 1520029804
transform 1 0 420 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1520029804
transform 1 0 404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1520029804
transform 1 0 428 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_135
timestamp 1520029804
transform 1 0 436 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_160
timestamp 1520029804
transform 1 0 444 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_138
timestamp 1520029804
transform 1 0 436 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1520029804
transform 1 0 460 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_174
timestamp 1520029804
transform 1 0 452 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_121
timestamp 1520029804
transform 1 0 484 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1520029804
transform 1 0 468 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1520029804
transform 1 0 476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1520029804
transform 1 0 532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1520029804
transform 1 0 548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1520029804
transform 1 0 540 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_139
timestamp 1520029804
transform 1 0 548 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1520029804
transform 1 0 540 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1520029804
transform 1 0 572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1520029804
transform 1 0 580 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_142
timestamp 1520029804
transform 1 0 580 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_143
timestamp 1520029804
transform 1 0 620 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1520029804
transform 1 0 628 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_128
timestamp 1520029804
transform 1 0 604 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_150
timestamp 1520029804
transform 1 0 612 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1520029804
transform 1 0 636 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_136
timestamp 1520029804
transform 1 0 612 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_163
timestamp 1520029804
transform 1 0 628 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_137
timestamp 1520029804
transform 1 0 636 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_180
timestamp 1520029804
transform 1 0 604 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_143
timestamp 1520029804
transform 1 0 628 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1520029804
transform 1 0 628 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1520029804
transform 1 0 660 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_181
timestamp 1520029804
transform 1 0 676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1520029804
transform 1 0 708 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1520029804
transform 1 0 740 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_146
timestamp 1520029804
transform 1 0 740 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1520029804
transform 1 0 772 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1520029804
transform 1 0 812 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1520029804
transform 1 0 764 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1520029804
transform 1 0 812 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_164
timestamp 1520029804
transform 1 0 772 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1520029804
transform 1 0 812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1520029804
transform 1 0 868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1520029804
transform 1 0 788 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_147
timestamp 1520029804
transform 1 0 812 0 1 385
box -3 -3 3 3
use turn_VIA0  turn_VIA0_8
timestamp 1520029804
transform 1 0 48 0 1 370
box -10 -3 10 3
use INVX2  INVX2_14
timestamp 1520029804
transform 1 0 72 0 1 370
box -9 -3 26 105
use NAND2X1  NAND2X1_0
timestamp 1520029804
transform -1 0 112 0 1 370
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_8
timestamp 1520029804
transform 1 0 112 0 1 370
box -8 -3 104 105
use FILL  FILL_62
timestamp 1520029804
transform 1 0 208 0 1 370
box -8 -3 16 105
use FILL  FILL_63
timestamp 1520029804
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_64
timestamp 1520029804
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_65
timestamp 1520029804
transform 1 0 232 0 1 370
box -8 -3 16 105
use FILL  FILL_66
timestamp 1520029804
transform 1 0 240 0 1 370
box -8 -3 16 105
use FILL  FILL_67
timestamp 1520029804
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_68
timestamp 1520029804
transform 1 0 256 0 1 370
box -8 -3 16 105
use FILL  FILL_69
timestamp 1520029804
transform 1 0 264 0 1 370
box -8 -3 16 105
use FILL  FILL_71
timestamp 1520029804
transform 1 0 272 0 1 370
box -8 -3 16 105
use FILL  FILL_72
timestamp 1520029804
transform 1 0 280 0 1 370
box -8 -3 16 105
use FILL  FILL_73
timestamp 1520029804
transform 1 0 288 0 1 370
box -8 -3 16 105
use INVX2  INVX2_15
timestamp 1520029804
transform 1 0 296 0 1 370
box -9 -3 26 105
use OAI21X1  OAI21X1_11
timestamp 1520029804
transform 1 0 312 0 1 370
box -8 -3 34 105
use INVX2  INVX2_16
timestamp 1520029804
transform 1 0 344 0 1 370
box -9 -3 26 105
use NAND3X1  NAND3X1_4
timestamp 1520029804
transform 1 0 360 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1520029804
transform 1 0 392 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_0
timestamp 1520029804
transform -1 0 456 0 1 370
box -8 -3 40 105
use M3_M2  M3_M2_148
timestamp 1520029804
transform 1 0 468 0 1 375
box -3 -3 3 3
use FILL  FILL_74
timestamp 1520029804
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_75
timestamp 1520029804
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_78
timestamp 1520029804
transform 1 0 472 0 1 370
box -8 -3 16 105
use FILL  FILL_80
timestamp 1520029804
transform 1 0 480 0 1 370
box -8 -3 16 105
use FILL  FILL_82
timestamp 1520029804
transform 1 0 488 0 1 370
box -8 -3 16 105
use FILL  FILL_84
timestamp 1520029804
transform 1 0 496 0 1 370
box -8 -3 16 105
use FILL  FILL_85
timestamp 1520029804
transform 1 0 504 0 1 370
box -8 -3 16 105
use INVX2  INVX2_17
timestamp 1520029804
transform 1 0 512 0 1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_8
timestamp 1520029804
transform -1 0 552 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1520029804
transform -1 0 576 0 1 370
box -8 -3 32 105
use M3_M2  M3_M2_149
timestamp 1520029804
transform 1 0 596 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_13
timestamp 1520029804
transform 1 0 576 0 1 370
box -8 -3 34 105
use NAND3X1  NAND3X1_7
timestamp 1520029804
transform -1 0 640 0 1 370
box -8 -3 40 105
use FILL  FILL_86
timestamp 1520029804
transform 1 0 640 0 1 370
box -8 -3 16 105
use FILL  FILL_87
timestamp 1520029804
transform 1 0 648 0 1 370
box -8 -3 16 105
use FILL  FILL_88
timestamp 1520029804
transform 1 0 656 0 1 370
box -8 -3 16 105
use FILL  FILL_89
timestamp 1520029804
transform 1 0 664 0 1 370
box -8 -3 16 105
use FILL  FILL_90
timestamp 1520029804
transform 1 0 672 0 1 370
box -8 -3 16 105
use FILL  FILL_91
timestamp 1520029804
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_92
timestamp 1520029804
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_93
timestamp 1520029804
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_94
timestamp 1520029804
transform 1 0 704 0 1 370
box -8 -3 16 105
use FILL  FILL_95
timestamp 1520029804
transform 1 0 712 0 1 370
box -8 -3 16 105
use FILL  FILL_96
timestamp 1520029804
transform 1 0 720 0 1 370
box -8 -3 16 105
use FILL  FILL_97
timestamp 1520029804
transform 1 0 728 0 1 370
box -8 -3 16 105
use FILL  FILL_98
timestamp 1520029804
transform 1 0 736 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_150
timestamp 1520029804
transform 1 0 756 0 1 375
box -3 -3 3 3
use FILL  FILL_99
timestamp 1520029804
transform 1 0 744 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_9
timestamp 1520029804
transform 1 0 752 0 1 370
box -8 -3 32 105
use M3_M2  M3_M2_151
timestamp 1520029804
transform 1 0 788 0 1 375
box -3 -3 3 3
use DFFPOSX1  DFFPOSX1_12
timestamp 1520029804
transform 1 0 776 0 1 370
box -8 -3 104 105
use FILL  FILL_100
timestamp 1520029804
transform 1 0 872 0 1 370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1520029804
transform 1 0 880 0 1 370
box -8 -3 16 105
use FILL  FILL_104
timestamp 1520029804
transform 1 0 888 0 1 370
box -8 -3 16 105
use turn_VIA0  turn_VIA0_9
timestamp 1520029804
transform 1 0 920 0 1 370
box -10 -3 10 3
use M3_M2  M3_M2_158
timestamp 1520029804
transform 1 0 76 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1520029804
transform 1 0 124 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1520029804
transform 1 0 84 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_160
timestamp 1520029804
transform 1 0 180 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1520029804
transform 1 0 204 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1520029804
transform 1 0 260 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_191
timestamp 1520029804
transform 1 0 180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1520029804
transform 1 0 108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1520029804
transform 1 0 164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1520029804
transform 1 0 204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1520029804
transform 1 0 260 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_152
timestamp 1520029804
transform 1 0 420 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1520029804
transform 1 0 388 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1520029804
transform 1 0 412 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1520029804
transform 1 0 380 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_192
timestamp 1520029804
transform 1 0 364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1520029804
transform 1 0 380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1520029804
transform 1 0 284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1520029804
transform 1 0 340 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_177
timestamp 1520029804
transform 1 0 388 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_215
timestamp 1520029804
transform 1 0 388 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_153
timestamp 1520029804
transform 1 0 444 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_185
timestamp 1520029804
transform 1 0 428 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1520029804
transform 1 0 412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1520029804
transform 1 0 428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1520029804
transform 1 0 412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1520029804
transform 1 0 404 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_183
timestamp 1520029804
transform 1 0 420 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_217
timestamp 1520029804
transform 1 0 444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1520029804
transform 1 0 436 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_164
timestamp 1520029804
transform 1 0 476 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_186
timestamp 1520029804
transform 1 0 476 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_178
timestamp 1520029804
transform 1 0 468 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_218
timestamp 1520029804
transform 1 0 468 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1520029804
transform 1 0 460 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1520029804
transform 1 0 452 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_154
timestamp 1520029804
transform 1 0 492 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1520029804
transform 1 0 484 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1520029804
transform 1 0 532 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1520029804
transform 1 0 524 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1520029804
transform 1 0 564 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_196
timestamp 1520029804
transform 1 0 532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1520029804
transform 1 0 556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1520029804
transform 1 0 564 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1520029804
transform 1 0 532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1520029804
transform 1 0 548 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_185
timestamp 1520029804
transform 1 0 524 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1520029804
transform 1 0 556 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1520029804
transform 1 0 588 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_199
timestamp 1520029804
transform 1 0 588 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1520029804
transform 1 0 580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1520029804
transform 1 0 596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1520029804
transform 1 0 540 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_186
timestamp 1520029804
transform 1 0 548 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1520029804
transform 1 0 612 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_187
timestamp 1520029804
transform 1 0 612 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1520029804
transform 1 0 644 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1520029804
transform 1 0 628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1520029804
transform 1 0 644 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_182
timestamp 1520029804
transform 1 0 628 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_223
timestamp 1520029804
transform 1 0 652 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_189
timestamp 1520029804
transform 1 0 652 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1520029804
transform 1 0 668 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_202
timestamp 1520029804
transform 1 0 668 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_155
timestamp 1520029804
transform 1 0 700 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1520029804
transform 1 0 716 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_203
timestamp 1520029804
transform 1 0 700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1520029804
transform 1 0 660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1520029804
transform 1 0 668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1520029804
transform 1 0 692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1520029804
transform 1 0 716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1520029804
transform 1 0 700 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_190
timestamp 1520029804
transform 1 0 700 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1520029804
transform 1 0 748 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1520029804
transform 1 0 740 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1520029804
transform 1 0 764 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_189
timestamp 1520029804
transform 1 0 748 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1520029804
transform 1 0 740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1520029804
transform 1 0 764 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1520029804
transform 1 0 740 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_180
timestamp 1520029804
transform 1 0 796 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1520029804
transform 1 0 828 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_206
timestamp 1520029804
transform 1 0 804 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1520029804
transform 1 0 820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1520029804
transform 1 0 780 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1520029804
transform 1 0 788 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_187
timestamp 1520029804
transform 1 0 788 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_231
timestamp 1520029804
transform 1 0 812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1520029804
transform 1 0 804 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_191
timestamp 1520029804
transform 1 0 780 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1520029804
transform 1 0 844 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_208
timestamp 1520029804
transform 1 0 844 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_176
timestamp 1520029804
transform 1 0 876 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_232
timestamp 1520029804
transform 1 0 860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1520029804
transform 1 0 852 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_188
timestamp 1520029804
transform 1 0 860 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_240
timestamp 1520029804
transform 1 0 876 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_192
timestamp 1520029804
transform 1 0 852 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_242
timestamp 1520029804
transform 1 0 868 0 1 305
box -2 -2 2 2
use turn_VIA0  turn_VIA0_10
timestamp 1520029804
transform 1 0 24 0 1 270
box -10 -3 10 3
use DFFPOSX1  DFFPOSX1_9
timestamp 1520029804
transform 1 0 72 0 -1 370
box -8 -3 104 105
use DFFPOSX1  DFFPOSX1_10
timestamp 1520029804
transform 1 0 168 0 -1 370
box -8 -3 104 105
use FILL  FILL_70
timestamp 1520029804
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_76
timestamp 1520029804
transform 1 0 272 0 -1 370
box -8 -3 16 105
use DFFPOSX1  DFFPOSX1_11
timestamp 1520029804
transform -1 0 376 0 -1 370
box -8 -3 104 105
use OAI21X1  OAI21X1_12
timestamp 1520029804
transform 1 0 376 0 -1 370
box -8 -3 34 105
use NOR2X1  NOR2X1_7
timestamp 1520029804
transform -1 0 432 0 -1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_6
timestamp 1520029804
transform 1 0 432 0 -1 370
box -8 -3 40 105
use FILL  FILL_77
timestamp 1520029804
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_79
timestamp 1520029804
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_81
timestamp 1520029804
transform 1 0 480 0 -1 370
box -8 -3 16 105
use FILL  FILL_83
timestamp 1520029804
transform 1 0 488 0 -1 370
box -8 -3 16 105
use FILL  FILL_102
timestamp 1520029804
transform 1 0 496 0 -1 370
box -8 -3 16 105
use AOI21X1  AOI21X1_2
timestamp 1520029804
transform -1 0 536 0 -1 370
box -7 -3 39 105
use NAND2X1  NAND2X1_2
timestamp 1520029804
transform -1 0 560 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_14
timestamp 1520029804
transform -1 0 592 0 -1 370
box -8 -3 34 105
use NOR2X1  NOR2X1_10
timestamp 1520029804
transform -1 0 616 0 -1 370
box -8 -3 32 105
use AOI21X1  AOI21X1_3
timestamp 1520029804
transform 1 0 616 0 -1 370
box -7 -3 39 105
use INVX2  INVX2_18
timestamp 1520029804
transform 1 0 648 0 -1 370
box -9 -3 26 105
use AOI21X1  AOI21X1_4
timestamp 1520029804
transform 1 0 664 0 -1 370
box -7 -3 39 105
use OAI21X1  OAI21X1_15
timestamp 1520029804
transform -1 0 728 0 -1 370
box -8 -3 34 105
use INVX2  INVX2_19
timestamp 1520029804
transform -1 0 744 0 -1 370
box -9 -3 26 105
use AOI21X1  AOI21X1_5
timestamp 1520029804
transform -1 0 776 0 -1 370
box -7 -3 39 105
use OAI21X1  OAI21X1_16
timestamp 1520029804
transform 1 0 776 0 -1 370
box -8 -3 34 105
use NOR2X1  NOR2X1_11
timestamp 1520029804
transform -1 0 832 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_20
timestamp 1520029804
transform -1 0 848 0 -1 370
box -9 -3 26 105
use NAND3X1  NAND3X1_8
timestamp 1520029804
transform 1 0 848 0 -1 370
box -8 -3 40 105
use FILL  FILL_103
timestamp 1520029804
transform 1 0 880 0 -1 370
box -8 -3 16 105
use FILL  FILL_105
timestamp 1520029804
transform 1 0 888 0 -1 370
box -8 -3 16 105
use turn_VIA0  turn_VIA0_11
timestamp 1520029804
transform 1 0 944 0 1 270
box -10 -3 10 3
use M2_M1  M2_M1_243
timestamp 1520029804
transform 1 0 124 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1520029804
transform 1 0 108 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1520029804
transform 1 0 100 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_215
timestamp 1520029804
transform 1 0 100 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_250
timestamp 1520029804
transform 1 0 140 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_203
timestamp 1520029804
transform 1 0 140 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_251
timestamp 1520029804
transform 1 0 172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1520029804
transform 1 0 148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1520029804
transform 1 0 156 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_204
timestamp 1520029804
transform 1 0 164 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_289
timestamp 1520029804
transform 1 0 156 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_216
timestamp 1520029804
transform 1 0 156 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_244
timestamp 1520029804
transform 1 0 204 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1520029804
transform 1 0 188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1520029804
transform 1 0 180 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_217
timestamp 1520029804
transform 1 0 188 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_252
timestamp 1520029804
transform 1 0 220 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_193
timestamp 1520029804
transform 1 0 316 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1520029804
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1520029804
transform 1 0 228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1520029804
transform 1 0 244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1520029804
transform 1 0 332 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_207
timestamp 1520029804
transform 1 0 284 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1520029804
transform 1 0 244 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1520029804
transform 1 0 316 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1520029804
transform 1 0 364 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_245
timestamp 1520029804
transform 1 0 348 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1520029804
transform 1 0 380 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1520029804
transform 1 0 348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1520029804
transform 1 0 364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1520029804
transform 1 0 372 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_198
timestamp 1520029804
transform 1 0 380 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_257
timestamp 1520029804
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1520029804
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1520029804
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1520029804
transform 1 0 372 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_208
timestamp 1520029804
transform 1 0 348 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1520029804
transform 1 0 396 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_259
timestamp 1520029804
transform 1 0 436 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_199
timestamp 1520029804
transform 1 0 444 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_277
timestamp 1520029804
transform 1 0 420 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_205
timestamp 1520029804
transform 1 0 436 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_278
timestamp 1520029804
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1520029804
transform 1 0 436 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_221
timestamp 1520029804
transform 1 0 436 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_260
timestamp 1520029804
transform 1 0 452 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_206
timestamp 1520029804
transform 1 0 460 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_261
timestamp 1520029804
transform 1 0 500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1520029804
transform 1 0 492 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_209
timestamp 1520029804
transform 1 0 492 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1520029804
transform 1 0 500 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1520029804
transform 1 0 556 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_247
timestamp 1520029804
transform 1 0 524 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1520029804
transform 1 0 524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1520029804
transform 1 0 532 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_210
timestamp 1520029804
transform 1 0 524 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_263
timestamp 1520029804
transform 1 0 596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1520029804
transform 1 0 660 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_200
timestamp 1520029804
transform 1 0 660 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_281
timestamp 1520029804
transform 1 0 556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1520029804
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1520029804
transform 1 0 660 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_211
timestamp 1520029804
transform 1 0 596 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1520029804
transform 1 0 532 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1520029804
transform 1 0 556 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1520029804
transform 1 0 620 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1520029804
transform 1 0 660 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_264
timestamp 1520029804
transform 1 0 692 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_201
timestamp 1520029804
transform 1 0 700 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_284
timestamp 1520029804
transform 1 0 700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1520029804
transform 1 0 764 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_196
timestamp 1520029804
transform 1 0 780 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_265
timestamp 1520029804
transform 1 0 740 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_202
timestamp 1520029804
transform 1 0 764 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1520029804
transform 1 0 876 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_266
timestamp 1520029804
transform 1 0 820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1520029804
transform 1 0 876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1520029804
transform 1 0 764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1520029804
transform 1 0 780 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1520029804
transform 1 0 796 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_213
timestamp 1520029804
transform 1 0 764 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1520029804
transform 1 0 756 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1520029804
transform 1 0 820 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1520029804
transform 1 0 796 0 1 185
box -3 -3 3 3
use turn_VIA0  turn_VIA0_12
timestamp 1520029804
transform 1 0 48 0 1 170
box -10 -3 10 3
use FILL  FILL_106
timestamp 1520029804
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_108
timestamp 1520029804
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_109
timestamp 1520029804
transform 1 0 88 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1520029804
transform 1 0 96 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_17
timestamp 1520029804
transform -1 0 152 0 1 170
box -8 -3 34 105
use NOR2X1  NOR2X1_13
timestamp 1520029804
transform 1 0 152 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1520029804
transform 1 0 176 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_18
timestamp 1520029804
transform -1 0 232 0 1 170
box -8 -3 34 105
use DFFPOSX1  DFFPOSX1_13
timestamp 1520029804
transform 1 0 232 0 1 170
box -8 -3 104 105
use INVX2  INVX2_21
timestamp 1520029804
transform 1 0 328 0 1 170
box -9 -3 26 105
use OAI21X1  OAI21X1_19
timestamp 1520029804
transform -1 0 376 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1520029804
transform -1 0 408 0 1 170
box -8 -3 34 105
use AOI21X1  AOI21X1_6
timestamp 1520029804
transform 1 0 408 0 1 170
box -7 -3 39 105
use INVX2  INVX2_22
timestamp 1520029804
transform 1 0 440 0 1 170
box -9 -3 26 105
use FILL  FILL_110
timestamp 1520029804
transform 1 0 456 0 1 170
box -8 -3 16 105
use FILL  FILL_119
timestamp 1520029804
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_121
timestamp 1520029804
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_123
timestamp 1520029804
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_124
timestamp 1520029804
transform 1 0 488 0 1 170
box -8 -3 16 105
use FILL  FILL_125
timestamp 1520029804
transform 1 0 496 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1520029804
transform 1 0 504 0 1 170
box -8 -3 32 105
use INVX2  INVX2_26
timestamp 1520029804
transform 1 0 528 0 1 170
box -9 -3 26 105
use DFFPOSX1  DFFPOSX1_15
timestamp 1520029804
transform 1 0 544 0 1 170
box -8 -3 104 105
use NAND2X1  NAND2X1_5
timestamp 1520029804
transform 1 0 640 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_24
timestamp 1520029804
transform -1 0 696 0 1 170
box -8 -3 34 105
use FILL  FILL_126
timestamp 1520029804
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_127
timestamp 1520029804
transform 1 0 704 0 1 170
box -8 -3 16 105
use FILL  FILL_128
timestamp 1520029804
transform 1 0 712 0 1 170
box -8 -3 16 105
use FILL  FILL_129
timestamp 1520029804
transform 1 0 720 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_25
timestamp 1520029804
transform 1 0 728 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_6
timestamp 1520029804
transform -1 0 784 0 1 170
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_16
timestamp 1520029804
transform 1 0 784 0 1 170
box -8 -3 104 105
use FILL  FILL_130
timestamp 1520029804
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_142
timestamp 1520029804
transform 1 0 888 0 1 170
box -8 -3 16 105
use turn_VIA0  turn_VIA0_13
timestamp 1520029804
transform 1 0 920 0 1 170
box -10 -3 10 3
use turn_VIA0  turn_VIA0_14
timestamp 1520029804
transform 1 0 24 0 1 70
box -10 -3 10 3
use M3_M2  M3_M2_231
timestamp 1520029804
transform 1 0 84 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_292
timestamp 1520029804
transform 1 0 84 0 1 135
box -2 -2 2 2
use FILL  FILL_107
timestamp 1520029804
transform 1 0 72 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_228
timestamp 1520029804
transform 1 0 132 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1520029804
transform 1 0 148 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1520029804
transform 1 0 140 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_293
timestamp 1520029804
transform 1 0 132 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1520029804
transform 1 0 140 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_294
timestamp 1520029804
transform 1 0 148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1520029804
transform 1 0 132 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1520029804
transform 1 0 140 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1520029804
transform 1 0 132 0 1 115
box -3 -3 3 3
use XNOR2X1  XNOR2X1_1
timestamp 1520029804
transform 1 0 80 0 -1 170
box -8 -3 64 105
use INVX2  INVX2_23
timestamp 1520029804
transform -1 0 152 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_230
timestamp 1520029804
transform 1 0 188 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1520029804
transform 1 0 196 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1520029804
transform 1 0 220 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_295
timestamp 1520029804
transform 1 0 180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1520029804
transform 1 0 188 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1520029804
transform 1 0 164 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1520029804
transform 1 0 180 0 1 105
box -3 -3 3 3
use OAI21X1  OAI21X1_21
timestamp 1520029804
transform 1 0 152 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_244
timestamp 1520029804
transform 1 0 204 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_297
timestamp 1520029804
transform 1 0 228 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1520029804
transform 1 0 236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1520029804
transform 1 0 212 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_252
timestamp 1520029804
transform 1 0 196 0 1 115
box -3 -3 3 3
use INVX2  INVX2_24
timestamp 1520029804
transform 1 0 184 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_312
timestamp 1520029804
transform 1 0 244 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_254
timestamp 1520029804
transform 1 0 236 0 1 105
box -3 -3 3 3
use OAI21X1  OAI21X1_22
timestamp 1520029804
transform 1 0 200 0 -1 170
box -8 -3 34 105
use INVX2  INVX2_25
timestamp 1520029804
transform 1 0 232 0 -1 170
box -9 -3 26 105
use FILL  FILL_111
timestamp 1520029804
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_112
timestamp 1520029804
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_113
timestamp 1520029804
transform 1 0 264 0 -1 170
box -8 -3 16 105
use FILL  FILL_114
timestamp 1520029804
transform 1 0 272 0 -1 170
box -8 -3 16 105
use FILL  FILL_115
timestamp 1520029804
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_116
timestamp 1520029804
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_117
timestamp 1520029804
transform 1 0 296 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_235
timestamp 1520029804
transform 1 0 356 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_299
timestamp 1520029804
transform 1 0 316 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1520029804
transform 1 0 420 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_300
timestamp 1520029804
transform 1 0 420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1520029804
transform 1 0 356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1520029804
transform 1 0 404 0 1 125
box -2 -2 2 2
use DFFPOSX1  DFFPOSX1_14
timestamp 1520029804
transform 1 0 304 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_245
timestamp 1520029804
transform 1 0 420 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_321
timestamp 1520029804
transform 1 0 420 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_3
timestamp 1520029804
transform 1 0 400 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_301
timestamp 1520029804
transform 1 0 452 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1520029804
transform 1 0 452 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_315
timestamp 1520029804
transform 1 0 460 0 1 125
box -2 -2 2 2
use OAI21X1  OAI21X1_23
timestamp 1520029804
transform -1 0 456 0 -1 170
box -8 -3 34 105
use FILL  FILL_118
timestamp 1520029804
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_120
timestamp 1520029804
transform 1 0 464 0 -1 170
box -8 -3 16 105
use FILL  FILL_122
timestamp 1520029804
transform 1 0 472 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_237
timestamp 1520029804
transform 1 0 516 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_302
timestamp 1520029804
transform 1 0 516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1520029804
transform 1 0 492 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_247
timestamp 1520029804
transform 1 0 516 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1520029804
transform 1 0 580 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1520029804
transform 1 0 620 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_303
timestamp 1520029804
transform 1 0 620 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1520029804
transform 1 0 540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1520029804
transform 1 0 580 0 1 125
box -2 -2 2 2
use OAI21X1  OAI21X1_26
timestamp 1520029804
transform 1 0 480 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_322
timestamp 1520029804
transform 1 0 516 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_7
timestamp 1520029804
transform -1 0 536 0 -1 170
box -8 -3 32 105
use DFFPOSX1  DFFPOSX1_17
timestamp 1520029804
transform -1 0 632 0 -1 170
box -8 -3 104 105
use FILL  FILL_131
timestamp 1520029804
transform 1 0 632 0 -1 170
box -8 -3 16 105
use FILL  FILL_132
timestamp 1520029804
transform 1 0 640 0 -1 170
box -8 -3 16 105
use FILL  FILL_133
timestamp 1520029804
transform 1 0 648 0 -1 170
box -8 -3 16 105
use FILL  FILL_134
timestamp 1520029804
transform 1 0 656 0 -1 170
box -8 -3 16 105
use FILL  FILL_135
timestamp 1520029804
transform 1 0 664 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_240
timestamp 1520029804
transform 1 0 684 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1520029804
transform 1 0 724 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_304
timestamp 1520029804
transform 1 0 684 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_248
timestamp 1520029804
transform 1 0 700 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1520029804
transform 1 0 788 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_305
timestamp 1520029804
transform 1 0 788 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1520029804
transform 1 0 724 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1520029804
transform 1 0 772 0 1 125
box -2 -2 2 2
use DFFPOSX1  DFFPOSX1_18
timestamp 1520029804
transform 1 0 672 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_249
timestamp 1520029804
transform 1 0 788 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_323
timestamp 1520029804
transform 1 0 788 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_8
timestamp 1520029804
transform 1 0 768 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_306
timestamp 1520029804
transform 1 0 820 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1520029804
transform 1 0 828 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_250
timestamp 1520029804
transform 1 0 820 0 1 125
box -3 -3 3 3
use OAI21X1  OAI21X1_27
timestamp 1520029804
transform -1 0 824 0 -1 170
box -8 -3 34 105
use INVX2  INVX2_27
timestamp 1520029804
transform 1 0 824 0 -1 170
box -9 -3 26 105
use FILL  FILL_136
timestamp 1520029804
transform 1 0 840 0 -1 170
box -8 -3 16 105
use FILL  FILL_137
timestamp 1520029804
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_138
timestamp 1520029804
transform 1 0 856 0 -1 170
box -8 -3 16 105
use FILL  FILL_139
timestamp 1520029804
transform 1 0 864 0 -1 170
box -8 -3 16 105
use FILL  FILL_140
timestamp 1520029804
transform 1 0 872 0 -1 170
box -8 -3 16 105
use FILL  FILL_141
timestamp 1520029804
transform 1 0 880 0 -1 170
box -8 -3 16 105
use FILL  FILL_143
timestamp 1520029804
transform 1 0 888 0 -1 170
box -8 -3 16 105
use turn_VIA0  turn_VIA0_15
timestamp 1520029804
transform 1 0 944 0 1 70
box -10 -3 10 3
use turn_VIA1  turn_VIA1_4
timestamp 1520029804
transform 1 0 48 0 1 47
box -10 -10 10 10
use turn_VIA1  turn_VIA1_5
timestamp 1520029804
transform 1 0 920 0 1 47
box -10 -10 10 10
use turn_VIA1  turn_VIA1_6
timestamp 1520029804
transform 1 0 24 0 1 23
box -10 -10 10 10
use turn_VIA1  turn_VIA1_7
timestamp 1520029804
transform 1 0 944 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal3 2 355 2 355 4 clka
rlabel metal2 116 838 116 838 4 clkb
rlabel metal3 2 405 2 405 4 restart
rlabel metal2 156 1 156 1 4 brake
rlabel metal2 140 1 140 1 4 left
rlabel metal2 180 1 180 1 4 right
rlabel metal2 332 1 332 1 4 l0
rlabel metal2 404 1 404 1 4 l1
rlabel metal2 540 1 540 1 4 l2
rlabel metal2 644 1 644 1 4 r0
rlabel metal3 966 215 966 215 4 r1
rlabel metal2 772 1 772 1 4 r2
rlabel metal2 564 838 564 838 4 error
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
<< end >>
